library ieee;
use ieee.std_logic_1164.all;

entity tb_xnor_gate is
end tb_xnor_gate;

architecture test of tb_xnor_gate is
	signal A,B,Y:std_logic;
	begin
		uut: entity work.xnor_gate
		port map(
			a=>A,
			b=>B,
			Y=>y
		);
		process
			begin
				A <= '0' ; B <= '0' ; wait for 10 ns;
				report "A = '0' , B = '0' , Y="&std_logic'image(Y);
				A <= '0' ; B <= '1' ; wait for 10 ns;
				report "A = '0' , B = '1' , Y="&std_logic'image(Y);
				A <= '1' ; B <= '0' ; wait for 10 ns;
				report "A = '1' , B = '0' , Y="&std_logic'image(Y);
				A <= '1' ; B <= '1' ; wait for 10 ns;
				report "A = '1' , B = '1' , Y="&std_logic'image(Y);
				wait;
		end process;
end architecture;