library ieee;
use ieee.std_logic_1164.all;

entity tb_xnor_gate is
end tb_xnor_gate;

architecture test of tb_xnor_gate is
	signal A,B,Y:std